module 7Seg_Decoder (
    input [3:0] sec_ones, sec_tens, mins,
    output [6:0] sec_ones_seg, sec_tens_seg, mins_seg
);

endmodule